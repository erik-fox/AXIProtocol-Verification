package axiprotocol;
  
class request;
	//What are the appropriate constraints
	rand bit [2:0] op;
	rand bit [31:0] address; 
	rand bit [3:0] readid;
	rand bit [3:0]readlen; 
	rand bit [2:0] readsize; 
	rand bit [1:0] readburst;
	rand bit [31:0]waddress; 
	rand bit [3:0] wlen;
	rand bit [3:0] wstrobe; 
	rand bit [2:0] wsize; 
	rand bit [1:0] wburst; 
	rand bit [31:0] data; 
	rand bit [3:0] writeid;
   // bit wlen_c[4] = '{2,4,8,16};
	//CONSTRAINTS
	//FROM THE SPEC:
	//AWLEN/ARLEN 0000 ->1 through 1111->16; wrapping bursts, length must be 2,4,8,16
	constraint AW_len{wlen dist {1:/11,2:/5, 3:/11, [4:6]:/15, 7:/11, [8:14]:/35, 15:/11 };}      //awlen 0001,0011,0111,1111
	constraint AR_len{readlen dist {1:/11,2:/5, 3:/11, [4:6]:/15, 7:/11,[8:14]:/35, 15:/11 };}   //arlen 0001,0011, 0111,1111
	//constraint Burst_len{wburst inside wlen_c;}											   //wrapping bursts, length must be 2,4,8,16
	//ARSIZE/AWSIZE 000->1 through 111 -> 128 size of transfer must not exceed data bus width in transaction
	constraint AR_size{readsize inside {[1:3]};}												//arsize 000, 001, 010
	constraint AW_size{wsize inside {[1:3]};}													//awsize 000, 001,010
	//ARBURST/AWBURST 00 -> fixed 01 -> INCR 10-> WRAP
	constraint AR_Burst{readburst inside {[0:2]};}												//arburst 00, 01, 10
	constraint AW_Burst{wburst inside {[0:2]};}													//awburst 00,01,10
	//IN THE CODE:
	//awaddr>32'h5ff and <=32'hfff and awsize <3'b100
	constraint AW_Addr{waddress inside {[32'h5ff:32'hfff]};}	
	//arsize 000, 001, 010
	//arburst 00, 01, 10
	//arlen 0001,0011, 0111,1111
	//awburst 00,01,10,
	//awsize 000, 001,010
	//awlen 0001,0011,0111,1111
	
	//araddr>32'h1ff aradddr<=32'hfff 
	constraint AR_Addr{address inside {[32'h1ff:32'hfff]};}
	//wstrb 0001, 0010, 0100,1000,0011,0101,1001, 0110, 1010,1100,00111,1110,1011, 1101, 1111,	
	constraint W_strobe{wstrobe inside {[1:15]};}
endclass// Code your design here
class tester;
	virtual tbbfm bfm;
    	function new(virtual tbbfm b);
      		bfm=b;
    	endfunction
	task execute();
		request r0;
		string testcase;

		r0=new();

		$value$plusargs("TESTCASE=%s",testcase);
		case(testcase)
			"readburst": read(32'h000005FF, 4'b0000, 4'b0000,3'b000,2'b00);//Read Burst 
			"overlapping_readburst":begin read(32'h000005FF, 4'b0000, 4'b0000,3'b000,2'b00);read(32'h00000600, 4'b0000, 4'b0000,3'b000,2'b00);end //overlapping readbursts
			"write_burst":write(32'h000006FE,4'b0011, 4'b0100, 3'b010,2'b01,32'hFFFFFFFF,4'b0100);//write burst
			"out_of_order":begin read(32'h000008FF, 4'b0001,4'b0011,3'b010,2'b01);write(32'h000006FE,4'b0011, 4'b0100, 3'b010,2'b01,32'hFFFFFFFF,4'b0100);end // Transaction ordering
			"fulltest":determine();
		endcase

		repeat(1000) 
		begin
          	@(posedge bfm.clk)
         	 begin
			assert(r0.randomize());
   
			case(r0.op)
				3'b000:read(r0.address,r0.readid, r0.readlen,r0.readsize,r0.readburst);//read
				3'b001: write(r0.waddress,r0.wlen, r0.wstrobe, r0.wsize,r0.wburst, r0.data, r0.writeid);//write
				3'b010: begin read(r0.address,r0.readid, r0.readlen,r0.readsize,r0.readburst);read(32'h00000600, 4'b0000, 4'b0000,3'b000,2'b00);end //overlapping readbursts
				3'b010: begin read(r0.address, r0.readid,r0.readlen,r0.readsize,r0.readburst);write(r0.waddress,r0.wlen, r0.wstrobe, r0.wsize,r0.wburst,r0.data,r0.writeid);end // Transaction ordering
			endcase
          	end
		end
	endtask
	task read(input bit [31:0] address, input bit[3:0] readid, input bit [3:0]readlen,input bit [2:0] readsize, input bit[1:0] readburst);
		@(negedge bfm.clk)begin
			bfm.araddr=address;
    			bfm.arid=readid;
    			bfm.arlen=readlen;
  			bfm.arsize=readsize;
  			bfm.arburst=readburst;
		end
	endtask
  
	task write(input bit [31:0]waddress, input bit [3:0] wlen, input bit [3:0] wstrobe, input bit [2:0] wsize, input bit [1:0] wburst, input bit [31:0] data, input bit [3:0] writeid);
		@(negedge bfm.clk)begin
			bfm.awaddr=waddress;
  			bfm.awlen=wlen;
	  		bfm.wstrb=wstrobe;
  			bfm.awsize=wsize;
			bfm.awburst=wburst;
 			bfm.wdata=data;
			bfm.awid=writeid;
		end
	endtask
	task determine();
		#50
		read(32'h00000FFF, 4'b0000, 4'b0000,3'b000,2'b00); //readburst
		#50
		read(32'h000005FF, 4'b0000, 4'b0000,3'b000,2'b00);//overlapping readburst
		read(32'h00000600, 4'b0000, 4'b0000,3'b000,2'b00);
		#50
		write(32'h000006FF,4'b0000, 4'b0000, 3'b000,2'b00,32'hFFFFFFFF,4'b0000);//write burst
    		#50	
		read(32'h000008FF, 4'b0000, 4'b0011,3'b000,2'b00);//variable read burst length
		#50
    		write(32'h000006FE,4'b0011, 4'b0000, 3'b000,2'b00,32'hFFFFFFFF,4'b0000);// variable write burst length
		#50
    		read(32'h000008FF, 4'b0000, 4'b0011,3'b000,2'b01);//variable read burst type
		#50
		write(32'h000006FE,4'b0011, 4'b0000, 3'b000,2'b01,32'hFFFFFFFF,4'b0000);// variable write burst type  
    		#50
		read(32'h000008FF, 4'b0000, 4'b0011,3'b010,2'b01);//variable read burst size
		#50
    		write(32'h000006FE,4'b0011, 4'b0000, 3'b010,2'b01,32'hFFFFFFFF,4'b0000);// variable write burst size
    		#50
    		read(32'h000008FF, 4'b0001,4'b0011,3'b010,2'b01);//Transaction ordering
	   	write(32'h000006FE,4'b0011, 4'b0100, 3'b010,2'b01,32'hFFFFFFFF,4'b0100);// Transaction ordering
		
		for(int i=32'h000006FF;i<=32'h00000FFF;i++) begin
			write(i,4'b0000, 4'b0000, 3'b000,2'b00,i,4'b0000);
		end
	
		#50
		read(32'h000006FF,4'b0000,4'b0100,3'b001,2'b00); //fixed read burst
		#50
		read(32'h000007FF,4'b0000,4'b0001,3'b000,2'b01); //incrementing read burst
		#50
		read(32'h00000700,4'b0000,4'b0001,3'b000,2'b10); //wrapping readburst
		//write and reading from same location
		#50
		write(32'h000006FF,4'b0000, 4'b0000, 3'b000,2'b00,32'hFFFFFFFF,4'b0000);
		read(32'h000006FF,4'b0000,4'b0000,3'b000,2'b00);
		//simultaneous write to different memory locations
		#50 
		write(32'h00000755,4'b0000, 4'b0000, 3'b000,2'b00,32'hFFFFFFFF,4'b0000);
		write(32'h00000765,4'b0000, 4'b0000, 3'b000,2'b00,32'hFFFFFFFF,4'b0000);
		//back to back writes to same memory and reading from it atlast
		#50 
		write(32'h000007EE,4'b0000, 4'b0000, 3'b000,2'b00,32'hFFF89000,4'b0000);
		write(32'h000007EE,4'b0000, 4'b0000, 3'b000,2'b00,32'hFFF89670,4'b0000);
		read(32'h000007EE,4'b0000,4'b0000,3'b000,2'b00);
		//Access out-of-bound memory
		#50
		read(32'hFFFFF7EE,4'b0000,4'b0000,3'b000,2'b00);
	endtask		
endclass 

class coverage;
	virtual tbbfm bfm;
	covergroup inputs;
		readaddr:coverpoint bfm.araddr;
		readid:coverpoint bfm.arid;
		readlen:coverpoint bfm.arlen;
		readsize:coverpoint bfm.arsize;
		readburst: coverpoint bfm.arburst;
		writeaddr:coverpoint bfm.awaddr;
		writelen:coverpoint bfm.awlen;
		writestrobe:coverpoint bfm.wstrb;
		writesize:coverpoint bfm.awsize;
		writeburst:coverpoint bfm.awburst;
		writedata:coverpoint bfm.wdata;
		writeid:coverpoint bfm.awid;
		read: cross readid, readlen, readsize, readburst;
		write: cross writelen, writestrobe, writesize, writeburst, writeid;
	endgroup
	covergroup outputs;
		//readburst
		readaddressvalid:coverpoint bfm.ARVALID;
		readaddressready:coverpoint bfm.ARREADY;
		readlast:coverpoint bfm.RLAST;
		readvalid:coverpoint bfm.RVALID;
		readready:coverpoint bfm.RREADY;
		readaddresssignals: cross readaddressvalid, readaddressready;
		readsignals: cross readvalid, readready;
		readsignalslast: cross readvalid, readready, readlast;
		//writeburst
		writeaddressvalid:coverpoint bfm.AWVALID;
		writeaddressready:coverpoint bfm.AWREADY;
		writelast: coverpoint bfm.WLAST;
		writevalid: coverpoint bfm.WVALID;
		writeready: coverpoint bfm.WREADY;
		writesignals: cross writevalid, writeready;
		writesignalslast: cross writelast, writevalid, writeready;
		writeresponse: coverpoint bfm.BRESP;
		writeresponsevalid: coverpoint bfm.BVALID;
		writeresponseready: coverpoint bfm.BREADY;
		writeresponsecross: cross writeresponse, writeresponsevalid, writeresponseready; 
	endgroup
	
	function new( virtual interface tbbfm b);
		inputs = new();
		outputs= new();
		bfm=b;
	endfunction
	task execute();
		forever begin
			@(posedge bfm.clk);
			inputs.sample();
			outputs.sample();
		end
	endtask 
endclass


class testbench;
	virtual tbbfm bfm;
	tester tester_h;
    	coverage coverage_h;
    	//scoreboard scoreboard_h;
	//checker checker_h;
    
    	function new (virtual tbbfm b);
      		bfm = b;
    	endfunction
    
    	task execute();
      		tester_h = new(bfm);
      		coverage_h= new(bfm);
      		//scoreboard_h = new(bfm);
		//checker_h = new(bfm);
      		fork
        		tester_h.execute();
        		coverage_h.execute();
        		//scoreboard_h.execute();
			//checker_h.execute();
      		join_none
    	endtask
endclass
  
	



endpackage
